----------------------------------------------------------------------------------
-- Company:        
-- Engineer:       simon.burkhardt
-- 
-- Create Date:    2023-04-21
-- Design Name:    skid buffer testbench
-- Module Name:    tb_axis - bh
-- Project Name:   
-- Target Devices: 
-- Tool Versions:  GHDL 0.37
-- Description:    
-- 
-- Dependencies:   
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

-- this testbench acts as a streaming master, sending bursts of data
-- counting from 1-4, also asserting tlast on the 4th data packet

-- the testbench itself acts as a correct streaming master which keeps the data
-- until it is acknowledged by the DUT by asserting tready.

-- the data pattern can be influenced by the user in 2 ways
-- + Tx requests are generated by changing the pattern in p_stimuli_tready
--   the master will try to send data for as long as sim_valid_data = '1'
-- + Rx acknowledgements are generated by changing the pattern in p_stimuli_tready
--   the downstream slave after the DUT will signal ready-to-receive 
--   when sim_ready_data = '1'

-- simulate both with OPT_DATA_REG = True / False
entity tb_axis is
  generic
  (
    OPT_DATA_REG         : boolean   := True;
    -- Width of ID for for write address, write data, read address and read data
    C_S_AXI_ID_WIDTH     : integer   := 3;
    -- Width of S_AXI data bus
    C_S_AXI_DATA_WIDTH   : integer   := 8;
    -- Width of S_AXI address bus
    C_S_AXI_ADDR_WIDTH   : integer   := 8;
    -- Width of optional user defined signal in write address channel
    C_S_AXI_AWUSER_WIDTH : integer   := 0;
    -- Width of optional user defined signal in read address channel
    C_S_AXI_ARUSER_WIDTH : integer   := 0;
    -- Width of optional user defined signal in write data channel
    C_S_AXI_WUSER_WIDTH  : integer   := 0;
    -- Width of optional user defined signal in read data channel
    C_S_AXI_RUSER_WIDTH  : integer   := 0;
    -- Width of optional user defined signal in write response channel
    C_S_AXI_BUSER_WIDTH  : integer   := 0
  );
end tb_axis;

architecture bh of tb_axis is
  -- DUT component declaration

  component axi4_s_write_splitter is
    generic (
      C_AXI_ID_WIDTH  : integer;
      C_AXI_DATA_WIDTH  : integer;
      C_AXI_ADDR_WIDTH  : integer;
      C_AXI_AWUSER_WIDTH  : integer;
      C_AXI_ARUSER_WIDTH  : integer;
      C_AXI_WUSER_WIDTH : integer;
      C_AXI_RUSER_WIDTH : integer;
      C_AXI_BUSER_WIDTH : integer
    );
    port (
      axi_aclk  : in std_logic;
      axi_aresetn : in std_logic;

      s00_axi_awid    : in std_logic_vector(C_AXI_ID_WIDTH-1 downto 0);
      s00_axi_awaddr  : in std_logic_vector(C_AXI_ADDR_WIDTH-1 downto 0);
      s00_axi_awlen   : in std_logic_vector(7 downto 0);
      s00_axi_awsize  : in std_logic_vector(2 downto 0);
      s00_axi_awburst : in std_logic_vector(1 downto 0);
      s00_axi_awlock  : in std_logic;
      s00_axi_awcache : in std_logic_vector(3 downto 0);
      s00_axi_awprot  : in std_logic_vector(2 downto 0);
      s00_axi_awqos   : in std_logic_vector(3 downto 0);
      s00_axi_awregion : in std_logic_vector(3 downto 0);
      s00_axi_awuser  : in std_logic_vector(C_AXI_AWUSER_WIDTH-1 downto 0);
      s00_axi_awvalid : in std_logic;
      s00_axi_awready : out std_logic;
      s00_axi_wdata   : in std_logic_vector(C_AXI_DATA_WIDTH-1 downto 0);
      s00_axi_wstrb   : in std_logic_vector((C_AXI_DATA_WIDTH/8)-1 downto 0);
      s00_axi_wlast   : in std_logic;
      s00_axi_wuser   : in std_logic_vector(C_AXI_WUSER_WIDTH-1 downto 0);
      s00_axi_wvalid  : in std_logic;
      s00_axi_wready  : out std_logic;
      s00_axi_bid     : out std_logic_vector(C_AXI_ID_WIDTH-1 downto 0);
      s00_axi_bresp   : out std_logic_vector(1 downto 0);
      s00_axi_buser   : out std_logic_vector(C_AXI_BUSER_WIDTH-1 downto 0);
      s00_axi_bvalid  : out std_logic;
      s00_axi_bready  : in std_logic;
      s00_axi_arid    : in std_logic_vector(C_AXI_ID_WIDTH-1 downto 0);
      s00_axi_araddr  : in std_logic_vector(C_AXI_ADDR_WIDTH-1 downto 0);
      s00_axi_arlen   : in std_logic_vector(7 downto 0);
      s00_axi_arsize  : in std_logic_vector(2 downto 0);
      s00_axi_arburst : in std_logic_vector(1 downto 0);
      s00_axi_arlock  : in std_logic;
      s00_axi_arcache : in std_logic_vector(3 downto 0);
      s00_axi_arprot  : in std_logic_vector(2 downto 0);
      s00_axi_arqos   : in std_logic_vector(3 downto 0);
      s00_axi_arregion : in std_logic_vector(3 downto 0);
      s00_axi_aruser  : in std_logic_vector(C_AXI_ARUSER_WIDTH-1 downto 0);
      s00_axi_arvalid : in std_logic;
      s00_axi_arready : out std_logic;
      s00_axi_rid     : out std_logic_vector(C_AXI_ID_WIDTH-1 downto 0);
      s00_axi_rdata   : out std_logic_vector(C_AXI_DATA_WIDTH-1 downto 0);
      s00_axi_rresp   : out std_logic_vector(1 downto 0);
      s00_axi_rlast   : out std_logic;
      s00_axi_ruser   : out std_logic_vector(C_AXI_RUSER_WIDTH-1 downto 0);
      s00_axi_rvalid  : out std_logic;
      s00_axi_rready  : in std_logic;
      
      m00_axi_awid    : out std_logic_vector(C_AXI_ID_WIDTH-1 downto 0);
      m00_axi_awaddr  : out std_logic_vector(C_AXI_ADDR_WIDTH-1 downto 0);
      m00_axi_awlen   : out std_logic_vector(7 downto 0);
      m00_axi_awsize  : out std_logic_vector(2 downto 0);
      m00_axi_awburst : out std_logic_vector(1 downto 0);
      m00_axi_awlock  : out std_logic;
      m00_axi_awcache : out std_logic_vector(3 downto 0);
      m00_axi_awprot  : out std_logic_vector(2 downto 0);
      m00_axi_awqos   : out std_logic_vector(3 downto 0);
      m00_axi_awuser  : out std_logic_vector(C_AXI_AWUSER_WIDTH-1 downto 0);
      m00_axi_awvalid : out std_logic;
      m00_axi_awready : in std_logic;
      m00_axi_wdata   : out std_logic_vector(C_AXI_DATA_WIDTH-1 downto 0);
      m00_axi_wstrb   : out std_logic_vector(C_AXI_DATA_WIDTH/8-1 downto 0);
      m00_axi_wlast   : out std_logic;
      m00_axi_wuser   : out std_logic_vector(C_AXI_WUSER_WIDTH-1 downto 0);
      m00_axi_wvalid  : out std_logic;
      m00_axi_wready  : in std_logic;
      m00_axi_bid     : in std_logic_vector(C_AXI_ID_WIDTH-1 downto 0);
      m00_axi_bresp   : in std_logic_vector(1 downto 0);
      m00_axi_buser   : in std_logic_vector(C_AXI_BUSER_WIDTH-1 downto 0);
      m00_axi_bvalid  : in std_logic;
      m00_axi_bready  : out std_logic;
      m00_axi_arid    : out std_logic_vector(C_AXI_ID_WIDTH-1 downto 0);
      m00_axi_araddr  : out std_logic_vector(C_AXI_ADDR_WIDTH-1 downto 0);
      m00_axi_arlen   : out std_logic_vector(7 downto 0);
      m00_axi_arsize  : out std_logic_vector(2 downto 0);
      m00_axi_arburst : out std_logic_vector(1 downto 0);
      m00_axi_arlock  : out std_logic;
      m00_axi_arcache : out std_logic_vector(3 downto 0);
      m00_axi_arprot  : out std_logic_vector(2 downto 0);
      m00_axi_arqos   : out std_logic_vector(3 downto 0);
      m00_axi_aruser  : out std_logic_vector(C_AXI_ARUSER_WIDTH-1 downto 0);
      m00_axi_arvalid : out std_logic;
      m00_axi_arready : in std_logic;
      m00_axi_rid     : in std_logic_vector(C_AXI_ID_WIDTH-1 downto 0);
      m00_axi_rdata   : in std_logic_vector(C_AXI_DATA_WIDTH-1 downto 0);
      m00_axi_rresp   : in std_logic_vector(1 downto 0);
      m00_axi_rlast   : in std_logic;
      m00_axi_ruser   : in std_logic_vector(C_AXI_RUSER_WIDTH-1 downto 0);
      m00_axi_rvalid  : in std_logic;
      m00_axi_rready  : out std_logic;

      m00_axis_tvalid : out std_logic;
      m00_axis_tdata  : out std_logic_vector(C_AXI_ADDR_WIDTH-1 downto 0);
      m00_axis_tstrb  : out std_logic_vector((C_AXI_ADDR_WIDTH/8)-1 downto 0);
      m00_axis_tlast  : out std_logic;
      m00_axis_tready : in std_logic;

      m01_axis_tvalid : out std_logic;
      m01_axis_tdata  : out std_logic_vector(C_AXI_DATA_WIDTH-1 downto 0);
      m01_axis_tstrb  : out std_logic_vector((C_AXI_DATA_WIDTH/8)-1 downto 0);
      m01_axis_tlast  : out std_logic;
      m01_axis_tready : in std_logic;

      m02_axis_tvalid : out std_logic;
      m02_axis_tdata  : out std_logic_vector(C_AXI_ADDR_WIDTH-1 downto 0);
      m02_axis_tstrb  : out std_logic_vector((C_AXI_ADDR_WIDTH/8)-1 downto 0);
      m02_axis_tlast  : out std_logic;
      m02_axis_tready : in std_logic;

      m03_axis_tvalid : out std_logic;
      m03_axis_tdata  : out std_logic_vector(C_AXI_DATA_WIDTH-1 downto 0);
      m03_axis_tstrb  : out std_logic_vector((C_AXI_DATA_WIDTH/8)-1 downto 0);
      m03_axis_tlast  : out std_logic;
      m03_axis_tready : in std_logic;

      opt_awready   : out std_logic;
      opt_wready    : out std_logic;
      opt_arready   : out std_logic;
      opt_rready    : out std_logic
    );
  end component;

  
  constant CLK_PERIOD: TIME := 5 ns;

  signal sim_start_write : std_logic := '0'; -- request AW channel
  signal sim_start_ready : std_logic := '0'; -- signal ready to receive from slave
  signal sim_valid_data  : std_logic := '0'; -- AW complete, now send W channel
  signal sim_data        : std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);

  signal o_axis_tvalid : std_logic;
  signal o_axis_tdata  : std_logic_vector(C_S_AXI_ADDR_WIDTH-1 downto 0);
  signal o_axis_tstrb  : std_logic_vector((C_S_AXI_ADDR_WIDTH/8)-1 downto 0);
  signal o_axis_tlast  : std_logic;
  signal i_axis_tready : std_logic := '0';

  signal clk   : std_logic;
  signal rst_n : std_logic;

  signal o_axi_awid     : std_logic_vector(C_S_AXI_ID_WIDTH-1 downto 0);
  signal o_axi_awaddr   : std_logic_vector(C_S_AXI_ADDR_WIDTH-1 downto 0);
  signal o_axi_awlen    : std_logic_vector(7 downto 0);
  signal o_axi_awsize   : std_logic_vector(2 downto 0);
  signal o_axi_awburst  : std_logic_vector(1 downto 0);
  signal o_axi_awlock   : std_logic;
  signal o_axi_awcache  : std_logic_vector(3 downto 0);
  signal o_axi_awprot   : std_logic_vector(2 downto 0);
  signal o_axi_awqos    : std_logic_vector(3 downto 0);
  signal o_axi_awregion : std_logic_vector(3 downto 0);
  signal o_axi_awuser   : std_logic_vector(C_S_AXI_AWUSER_WIDTH-1 downto 0);
  signal o_axi_awvalid  : std_logic;
  signal i_axi_awready  : std_logic;
  signal o_axi_wdata    : std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
  signal o_axi_wstrb    : std_logic_vector((C_S_AXI_DATA_WIDTH/8)-1 downto 0);
  signal o_axi_wlast    : std_logic;
  signal o_axi_wuser    : std_logic_vector(C_S_AXI_WUSER_WIDTH-1 downto 0);
  signal o_axi_wvalid   : std_logic;
  signal i_axi_wready   : std_logic;
  signal i_axi_bid      : std_logic_vector(C_S_AXI_ID_WIDTH-1 downto 0);
  signal i_axi_bresp    : std_logic_vector(1 downto 0);
  signal i_axi_buser    : std_logic_vector(C_S_AXI_BUSER_WIDTH-1 downto 0);
  signal i_axi_bvalid   : std_logic;
  signal o_axi_bready   : std_logic;
  signal o_axi_arid     : std_logic_vector(C_S_AXI_ID_WIDTH-1 downto 0);
  signal o_axi_araddr   : std_logic_vector(C_S_AXI_ADDR_WIDTH-1 downto 0);
  signal o_axi_arlen    : std_logic_vector(7 downto 0);
  signal o_axi_arsize   : std_logic_vector(2 downto 0);
  signal o_axi_arburst  : std_logic_vector(1 downto 0);
  signal o_axi_arlock   : std_logic;
  signal o_axi_arcache  : std_logic_vector(3 downto 0);
  signal o_axi_arprot   : std_logic_vector(2 downto 0);
  signal o_axi_arqos    : std_logic_vector(3 downto 0);
  signal o_axi_arregion : std_logic_vector(3 downto 0);
  signal o_axi_aruser   : std_logic_vector(C_S_AXI_ARUSER_WIDTH-1 downto 0);
  signal o_axi_arvalid  : std_logic;
  signal i_axi_arready  : std_logic;
  signal i_axi_rid      : std_logic_vector(C_S_AXI_ID_WIDTH-1 downto 0);
  signal i_axi_rdata    : std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
  signal i_axi_rresp    : std_logic_vector(1 downto 0);
  signal i_axi_rlast    : std_logic;
  signal i_axi_ruser    : std_logic_vector(C_S_AXI_RUSER_WIDTH-1 downto 0);
  signal i_axi_rvalid   : std_logic;
  signal o_axi_rready   : std_logic;

  signal o_Y_axi_awid     : std_logic_vector(C_S_AXI_ID_WIDTH-1 downto 0);
  signal o_Y_axi_awaddr   : std_logic_vector(C_S_AXI_ADDR_WIDTH-1 downto 0);
  signal o_Y_axi_awlen    : std_logic_vector(7 downto 0);
  signal o_Y_axi_awsize   : std_logic_vector(2 downto 0);
  signal o_Y_axi_awburst  : std_logic_vector(1 downto 0);
  signal o_Y_axi_awlock   : std_logic;
  signal o_Y_axi_awcache  : std_logic_vector(3 downto 0);
  signal o_Y_axi_awprot   : std_logic_vector(2 downto 0);
  signal o_Y_axi_awqos    : std_logic_vector(3 downto 0);
  signal o_Y_axi_awregion : std_logic_vector(3 downto 0);
  signal o_Y_axi_awuser   : std_logic_vector(C_S_AXI_AWUSER_WIDTH-1 downto 0);
  signal o_Y_axi_awvalid  : std_logic;
  signal i_Y_axi_awready  : std_logic;
  signal o_Y_axi_wdata    : std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
  signal o_Y_axi_wstrb    : std_logic_vector((C_S_AXI_DATA_WIDTH/8)-1 downto 0);
  signal o_Y_axi_wlast    : std_logic;
  signal o_Y_axi_wuser    : std_logic_vector(C_S_AXI_WUSER_WIDTH-1 downto 0);
  signal o_Y_axi_wvalid   : std_logic;
  signal i_Y_axi_wready   : std_logic;
  signal i_Y_axi_bid      : std_logic_vector(C_S_AXI_ID_WIDTH-1 downto 0);
  signal i_Y_axi_bresp    : std_logic_vector(1 downto 0);
  signal i_Y_axi_buser    : std_logic_vector(C_S_AXI_BUSER_WIDTH-1 downto 0);
  signal i_Y_axi_bvalid   : std_logic;
  signal o_Y_axi_bready   : std_logic;
  signal o_Y_axi_arid     : std_logic_vector(C_S_AXI_ID_WIDTH-1 downto 0);
  signal o_Y_axi_araddr   : std_logic_vector(C_S_AXI_ADDR_WIDTH-1 downto 0);
  signal o_Y_axi_arlen    : std_logic_vector(7 downto 0);
  signal o_Y_axi_arsize   : std_logic_vector(2 downto 0);
  signal o_Y_axi_arburst  : std_logic_vector(1 downto 0);
  signal o_Y_axi_arlock   : std_logic;
  signal o_Y_axi_arcache  : std_logic_vector(3 downto 0);
  signal o_Y_axi_arprot   : std_logic_vector(2 downto 0);
  signal o_Y_axi_arqos    : std_logic_vector(3 downto 0);
  signal o_Y_axi_arregion : std_logic_vector(3 downto 0);
  signal o_Y_axi_aruser   : std_logic_vector(C_S_AXI_ARUSER_WIDTH-1 downto 0);
  signal o_Y_axi_arvalid  : std_logic;
  signal i_Y_axi_arready  : std_logic;
  signal i_Y_axi_rid      : std_logic_vector(C_S_AXI_ID_WIDTH-1 downto 0);
  signal i_Y_axi_rdata    : std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
  signal i_Y_axi_rresp    : std_logic_vector(1 downto 0);
  signal i_Y_axi_rlast    : std_logic;
  signal i_Y_axi_ruser    : std_logic_vector(C_S_AXI_RUSER_WIDTH-1 downto 0);
  signal i_Y_axi_rvalid   : std_logic;
  signal o_Y_axi_rready   : std_logic;

  signal clk_count : std_logic_vector(7 downto 0) := (others => '0');
  signal outstanding_xfers : std_logic_vector(7 downto 0) := (others => '0');
begin

  -- generate clk signal
  p_clk_gen : process
  begin
   clk <= '1';
   wait for (CLK_PERIOD / 2);
   clk <= '0';
   wait for (CLK_PERIOD / 2);
   clk_count <= std_logic_vector(unsigned(clk_count) + 1);
  end process;

  -- generate initial reset
  p_reset_gen : process
  begin 
    rst_n <= '0';
    wait until rising_edge(clk);
    wait for (CLK_PERIOD / 4);
    rst_n <= '1';
    wait;
  end process;

  axi4_s_axis_s_splitter_inst : axi4_s_write_splitter
    generic map (
      C_AXI_ID_WIDTH      => C_S_AXI_ID_WIDTH, 
      C_AXI_DATA_WIDTH    => C_S_AXI_DATA_WIDTH, 
      C_AXI_ADDR_WIDTH    => C_S_AXI_ADDR_WIDTH, 
      C_AXI_AWUSER_WIDTH  => C_S_AXI_AWUSER_WIDTH, 
      C_AXI_ARUSER_WIDTH  => C_S_AXI_ARUSER_WIDTH, 
      C_AXI_WUSER_WIDTH   => C_S_AXI_WUSER_WIDTH, 
      C_AXI_RUSER_WIDTH   => C_S_AXI_RUSER_WIDTH, 
      C_AXI_BUSER_WIDTH   => C_S_AXI_BUSER_WIDTH
    )
    port map (
      axi_aclk    => clk,
      axi_aresetn => rst_n,

      s00_axi_awid      => (others => '0'), -- o_axi_awid,        --n std_logic_vector(C_AXI_ID_WIDTH-1 downto 0);
      s00_axi_awaddr    => (others => '0'), -- o_axi_awaddr,        --n std_logic_vector(C_AXI_ADDR_WIDTH-1 downto 0);
      s00_axi_awlen     => (others => '0'), -- o_axi_awlen,        --n std_logic_vector(7 downto 0);
      s00_axi_awsize    => (others => '0'), -- o_axi_awsize,        --n std_logic_vector(2 downto 0);
      s00_axi_awburst   => (others => '0'), -- o_axi_awburst,        --n std_logic_vector(1 downto 0);
      s00_axi_awlock    => '0', -- o_axi_awlock,        --n std_logic;
      s00_axi_awcache   => (others => '0'), -- o_axi_awcache,        --n std_logic_vector(3 downto 0);
      s00_axi_awprot    => (others => '0'), -- o_axi_awprot,        --n std_logic_vector(2 downto 0);
      s00_axi_awqos     => (others => '0'), -- o_axi_awqos,        --n std_logic_vector(3 downto 0);
      s00_axi_awregion  => (others => '0'), -- o_axi_awregion,        --n std_logic_vector(3 downto 0);
      s00_axi_awuser    => (others => '0'), -- o_axi_awuser,        --n std_logic_vector(C_AXI_AWUSER_WIDTH-1 downto 0);
      s00_axi_awvalid   => '0', -- o_axi_awvalid,        --n std_logic;
      s00_axi_awready   => open, -- i_axi_awready,        --ut std_logic;
      s00_axi_wdata     => (others => '0'), -- o_axi_wdata,        --n std_logic_vector(C_AXI_DATA_WIDTH-1 downto 0);
      s00_axi_wstrb     => (others => '0'), -- o_axi_wstrb,        --n std_logic_vector((C_AXI_DATA_WIDTH/8)-1 downto 0);
      s00_axi_wlast     => '0', -- o_axi_wlast,        --n std_logic;
      s00_axi_wuser     => (others => '0'), -- o_axi_wuser,        --n std_logic_vector(C_AXI_WUSER_WIDTH-1 downto 0);
      s00_axi_wvalid    => '0', -- o_axi_wvalid,        --n std_logic;
      s00_axi_wready    => open, -- i_axi_wready,        --ut std_logic;
      s00_axi_bid       => open, -- i_axi_bid,        --ut std_logic_vector(C_AXI_ID_WIDTH-1 downto 0);
      s00_axi_bresp     => open, -- i_axi_bresp,        --ut std_logic_vector(1 downto 0);
      s00_axi_buser     => open, -- i_axi_buser,        --ut std_logic_vector(C_AXI_BUSER_WIDTH-1 downto 0);
      s00_axi_bvalid    => open, -- i_axi_bvalid,        --ut std_logic;
      s00_axi_bready    => '0', -- o_axi_bready,        --n std_logic;
      s00_axi_arid      => (others => '0'), -- o_axi_arid,        --n std_logic_vector(C_AXI_ID_WIDTH-1 downto 0);
      s00_axi_araddr    => (others => '0'), -- o_axi_araddr,        --n std_logic_vector(C_AXI_ADDR_WIDTH-1 downto 0);
      s00_axi_arlen     => (others => '0'), -- o_axi_arlen,        --n std_logic_vector(7 downto 0);
      s00_axi_arsize    => (others => '0'), -- o_axi_arsize,        --n std_logic_vector(2 downto 0);
      s00_axi_arburst   => (others => '0'), -- o_axi_arburst,        --n std_logic_vector(1 downto 0);
      s00_axi_arlock    => '0', -- o_axi_arlock,        --n std_logic;
      s00_axi_arcache   => (others => '0'), -- o_axi_arcache,        --n std_logic_vector(3 downto 0);
      s00_axi_arprot    => (others => '0'), -- o_axi_arprot,        --n std_logic_vector(2 downto 0);
      s00_axi_arqos     => (others => '0'), -- o_axi_arqos,        --n std_logic_vector(3 downto 0);
      s00_axi_arregion  => (others => '0'), -- o_axi_arregion,        --n std_logic_vector(3 downto 0);
      s00_axi_aruser    => (others => '0'), -- o_axi_aruser,        --n std_logic_vector(C_AXI_ARUSER_WIDTH-1 downto 0);
      s00_axi_arvalid   => '0', -- o_axi_arvalid,        --n std_logic;
      s00_axi_arready   => open, -- i_axi_arready,        --ut std_logic;
      s00_axi_rid       => open, -- i_axi_rid,        --ut std_logic_vector(C_AXI_ID_WIDTH-1 downto 0);
      s00_axi_rdata     => open, -- i_axi_rdata,        --ut std_logic_vector(C_AXI_DATA_WIDTH-1 downto 0);
      s00_axi_rresp     => open, -- i_axi_rresp,        --ut std_logic_vector(1 downto 0);
      s00_axi_rlast     => open, -- i_axi_rlast,        --ut std_logic;
      s00_axi_ruser     => open, -- i_axi_ruser,        --ut std_logic_vector(C_AXI_RUSER_WIDTH-1 downto 0);
      s00_axi_rvalid    => open, -- i_axi_rvalid,        --ut std_logic;
      s00_axi_rready    => '0', -- o_axi_rready,        --n std_logic;
      
      m00_axi_awid    => open, -- o_Y_axi_awid, --         ut std_logic_vector(C_AXI_ID_WIDTH-1 downto 0);
      m00_axi_awaddr  => open, -- o_Y_axi_awaddr, --         ut std_logic_vector(C_AXI_ADDR_WIDTH-1 downto 0);
      m00_axi_awlen   => open, -- o_Y_axi_awlen, --         ut std_logic_vector(7 downto 0);
      m00_axi_awsize  => open, -- o_Y_axi_awsize, --         ut std_logic_vector(2 downto 0);
      m00_axi_awburst => open, -- o_Y_axi_awburst, --         ut std_logic_vector(1 downto 0);
      m00_axi_awlock  => open, -- o_Y_axi_awlock, --         ut std_logic;
      m00_axi_awcache => open, -- o_Y_axi_awcache, --         ut std_logic_vector(3 downto 0);
      m00_axi_awprot  => open, -- o_Y_axi_awprot, --         ut std_logic_vector(2 downto 0);
      m00_axi_awqos   => open, -- o_Y_axi_awqos, --         ut std_logic_vector(3 downto 0);
      m00_axi_awuser  => open, -- o_Y_axi_awuser, --         ut std_logic_vector(C_AXI_AWUSER_WIDTH-1 downto 0);
      m00_axi_awvalid => open, -- o_Y_axi_awvalid, --         ut std_logic;
      m00_axi_awready => '0', -- i_Y_axi_awready, --         n std_logic;
      m00_axi_wdata   => open, -- o_Y_axi_wdata, --         ut std_logic_vector(C_AXI_DATA_WIDTH-1 downto 0);
      m00_axi_wstrb   => open, -- o_Y_axi_wstrb, --         ut std_logic_vector(C_AXI_DATA_WIDTH/8-1 downto 0);
      m00_axi_wlast   => open, -- o_Y_axi_wlast, --         ut std_logic;
      m00_axi_wuser   => open, -- o_Y_axi_wuser, --         ut std_logic_vector(C_AXI_WUSER_WIDTH-1 downto 0);
      m00_axi_wvalid  => open, -- o_Y_axi_wvalid, --         ut std_logic;
      m00_axi_wready  => '0', -- i_Y_axi_wready, --         n std_logic;
      m00_axi_bid     => (others => '0'), -- i_Y_axi_bid, --         n std_logic_vector(C_AXI_ID_WIDTH-1 downto 0);
      m00_axi_bresp   => (others => '0'), -- i_Y_axi_bresp, --         n std_logic_vector(1 downto 0);
      m00_axi_buser   => (others => '0'), -- i_Y_axi_buser, --         n std_logic_vector(C_AXI_BUSER_WIDTH-1 downto 0);
      m00_axi_bvalid  => '0', -- i_Y_axi_bvalid, --         n std_logic;
      m00_axi_bready  => open, -- o_Y_axi_bready, --         ut std_logic;
      m00_axi_arid    => open, -- o_Y_axi_arid, --         ut std_logic_vector(C_AXI_ID_WIDTH-1 downto 0);
      m00_axi_araddr  => open, -- o_Y_axi_araddr, --         ut std_logic_vector(C_AXI_ADDR_WIDTH-1 downto 0);
      m00_axi_arlen   => open, -- o_Y_axi_arlen, --         ut std_logic_vector(7 downto 0);
      m00_axi_arsize  => open, -- o_Y_axi_arsize, --         ut std_logic_vector(2 downto 0);
      m00_axi_arburst => open, -- o_Y_axi_arburst, --         ut std_logic_vector(1 downto 0);
      m00_axi_arlock  => open, -- o_Y_axi_arlock, --         ut std_logic;
      m00_axi_arcache => open, -- o_Y_axi_arcache, --         ut std_logic_vector(3 downto 0);
      m00_axi_arprot  => open, -- o_Y_axi_arprot, --         ut std_logic_vector(2 downto 0);
      m00_axi_arqos   => open, -- o_Y_axi_arqos, --         ut std_logic_vector(3 downto 0);
      m00_axi_aruser  => open, -- o_Y_axi_aruser, --         ut std_logic_vector(C_AXI_ARUSER_WIDTH-1 downto 0);
      m00_axi_arvalid => open, -- o_Y_axi_arvalid, --         ut std_logic;
      m00_axi_arready => '0', -- i_Y_axi_arready, --         n std_logic;
      m00_axi_rid     => (others => '0'), -- i_Y_axi_rid, --         n std_logic_vector(C_AXI_ID_WIDTH-1 downto 0);
      m00_axi_rdata   => (others => '0'), -- i_Y_axi_rdata, --         n std_logic_vector(C_AXI_DATA_WIDTH-1 downto 0);
      m00_axi_rresp   => (others => '0'), -- i_Y_axi_rresp, --         n std_logic_vector(1 downto 0);
      m00_axi_rlast   => '0', -- i_Y_axi_rlast, --         n std_logic;
      m00_axi_ruser   => (others => '0'), -- i_Y_axi_ruser, --         n std_logic_vector(C_AXI_RUSER_WIDTH-1 downto 0);
      m00_axi_rvalid  => '0', -- i_Y_axi_rvalid, --         n std_logic;
      m00_axi_rready  => open, -- o_Y_axi_rready, --         ut std_logic;

      m00_axis_tvalid => open, -- ;
      m00_axis_tdata  => open, -- (C_AXI_ADDR_WIDTH-1 downto 0);
      m00_axis_tstrb  => open, -- ((C_AXI_ADDR_WIDTH/8)-1 downto 0);
      m00_axis_tlast  => open, -- ;
      m00_axis_tready => '1',

      m01_axis_tvalid => open, -- ;
      m01_axis_tdata  => open, -- (C_AXI_DATA_WIDTH-1 downto 0);
      m01_axis_tstrb  => open, -- ((C_AXI_DATA_WIDTH/8)-1 downto 0);
      m01_axis_tlast  => open, -- ;
      m01_axis_tready => '1',

      m02_axis_tvalid => open, -- ;
      m02_axis_tdata  => open, -- (C_AXI_ADDR_WIDTH-1 downto 0);
      m02_axis_tstrb  => open, -- ((C_AXI_ADDR_WIDTH/8)-1 downto 0);
      m02_axis_tlast  => open, -- ;
      m02_axis_tready => '1',

      m03_axis_tvalid => open, -- ;
      m03_axis_tdata  => open, -- (C_AXI_DATA_WIDTH-1 downto 0);
      m03_axis_tstrb  => open, -- ((C_AXI_DATA_WIDTH/8)-1 downto 0);
      m03_axis_tlast  => open, -- ;
      m03_axis_tready => '1',

      opt_awready   => open,
      opt_wready    => open,
      opt_arready   => open,
      opt_rready    => open
    );
    
end bh;
